module sprites(
	input logic [5:0]          n_sprite,
	input logic [9:0]          line,
	input logic                clk,
	output logic [31:0][23:0]  pattern);

	always_ff @(posedge clk) begin
		case (n_sprite)
			6'd1 : begin
				case(line)
					10'd0 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h2d2d06}, {24'h605f06}, {24'h646305}, {24'h595806}, {24'h3e3d07}, {24'h090903}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd1 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h050506}, {24'h58666c}, {24'hcbd54f}, {24'hfdfc06}, {24'hfffd00}, {24'hfffd02}, {24'hf4f203}, {24'hd1cf07}, {24'h5f5e07}, {24'h000000}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd2 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h536375}, {24'hb2d6fe}, {24'hb3d6fb}, {24'hcde3a7}, {24'hfefd04}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfaf801}, {24'h686709}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd3 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h1f252b}, {24'ha4c5e9}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hd8e984}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hf1ef03}, {24'h2d2d05}, {24'h000000}, {10{24'h0}}};
					10'd4 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h66798f}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hb2d6fe}, {24'ha6c7ea}, {24'h242403}, {24'ha09f01}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'h818007}, {24'h000000}, {10{24'h0}}};
					10'd5 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h88a3c0}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hb4d7f8}, {24'hb9d3bd}, {24'h474702}, {24'hafad00}, {24'hfffd00}, {24'hfffd00}, {24'hfde937}, {24'hc59f79}, {24'h181215}, {10{24'h0}}};
					10'd6 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h8eaac9}, {24'hb2d6fe}, {24'hb2d6fe}, {24'hbddcda}, {24'hedf43b}, {24'hfefc05}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfef220}, {24'hf6b2d1}, {24'hf6b0d6}, {24'h664a5a}, {10{24'h0}}};
					10'd7 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h020202}, {24'h96b3d4}, {24'hb2d6fe}, {24'hcde4a6}, {24'hf9fa14}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfad56f}, {24'hf6b0d6}, {24'hf6b0d6}, {24'h8a6479}, {10{24'h0}}};
					10'd8 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h070809}, {24'h9bbadd}, {24'hbadae4}, {24'hfafb10}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfacd85}, {24'hf6b0d6}, {24'hf6b0d6}, {24'h9a6f87}, {10{24'h0}}};
					10'd9 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h070809}, {24'h9fbcd0}, {24'he4ef5a}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfdf21f}, {24'hca92af}, {24'hf6b0d6}, {24'h966d83}, {10{24'h0}}};
					10'd10 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h040404}, {24'hbbc868}, {24'hfffd01}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hf8f707}, {24'h31252b}, {24'he9a7ca}, {24'h775769}, {10{24'h0}}};
					10'd11 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h1c1c03}, {24'hf1ef03}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd03}, {24'h20200b}, {24'h7a596b}, {24'h21181d}, {10{24'h0}}};
					10'd12 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h3a3905}, {24'hfefc01}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd01}, {24'hfffd00}, {24'hfffd00}, {24'hfffd05}, {24'h636218}, {24'h030203}, {24'h000000}, {10{24'h0}}};
					10'd13 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h99980a}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd00}, {24'hfffd24}, {24'hfefd86}, {24'hb2b17c}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd14 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h1a1a06}, {24'hfcfa03}, {24'hfffd00}, {24'hfffd00}, {24'hfefd53}, {24'hfefd6e}, {24'hfffd6d}, {24'hfefd72}, {24'hfefd80}, {24'hfefd96}, {24'hfefdb1}, {24'hfefdb2}, {24'hf3f2ab}, {24'h222219}, {24'h000000}, {10{24'h0}}};
					10'd15 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h555407}, {24'hfffd00}, {24'hfffd00}, {24'hfffd28}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'h57573e}, {24'h000000}, {10{24'h0}}};
					10'd16 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h949308}, {24'hfffd00}, {24'hfffd08}, {24'hfefd7b}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd75}, {24'hfefd7b}, {24'hfefdb1}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'h83835d}, {24'h000000}, {10{24'h0}}};
					10'd17 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'hd7d608}, {24'hfffd00}, {24'hfffd39}, {24'hfefdb1}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfffd3c}, {24'hfffd06}, {24'hfdfc66}, {24'hfdfdb3}, {24'hfefdb2}, {24'hfefdb2}, {24'hbbba84}, {24'h000000}, {10{24'h0}}};
					10'd18 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h1a1a06}, {24'hfffd01}, {24'hfffd05}, {24'hfefd8a}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd6d}, {24'hfffd00}, {24'hedf43c}, {24'hbedcef}, {24'hf9fbb7}, {24'hfefdb2}, {24'hdfde9d}, {24'h161611}, {10{24'h0}}};
					10'd19 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h525209}, {24'hfffd00}, {24'hfffd28}, {24'hfefdb0}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd89}, {24'hfffd00}, {24'hf8f918}, {24'hb8d9ec}, {24'hdcecd4}, {24'hfefdb2}, {24'hebeaa5}, {24'h2e2e22}, {10{24'h0}}};
					10'd20 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h7b7a09}, {24'hfffd00}, {24'hfffd66}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd8a}, {24'hfffd00}, {24'hf9fa15}, {24'hb9dae7}, {24'hdfedd2}, {24'hfefdb2}, {24'hebeba6}, {24'h2f2e22}, {10{24'h0}}};
					10'd21 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'haeac0b}, {24'hfffd07}, {24'hfefda6}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb1}, {24'hfefd72}, {24'hfffd00}, {24'hf6f91e}, {24'hb6d8f1}, {24'heff5be}, {24'hfefdb2}, {24'hdede9d}, {24'h151510}, {10{24'h0}}};
					10'd22 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'hc8c707}, {24'hfffd20}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb1}, {24'hfffd29}, {24'hfffd00}, {24'he0ed67}, {24'hbddbf0}, {24'hfefdb1}, {24'hfefdb2}, {24'hcccc91}, {24'h000000}, {10{24'h0}}};
					10'd23 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h0b0a03}, {24'hdfdd04}, {24'hfefd33}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd7e}, {24'hfffd02}, {24'hfafb10}, {24'hc0ddd5}, {24'he6f1c9}, {24'hfefdb2}, {24'hfefdb2}, {24'hbfbe87}, {24'h000000}, {10{24'h0}}};
					10'd24 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h212103}, {24'hf6f407}, {24'hfefd58}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefda9}, {24'hfffd1c}, {24'hfffd00}, {24'hd5e88b}, {24'hcde4e1}, {24'hfdfdb3}, {24'hfefdb2}, {24'hfefdb2}, {24'hb4b37f}, {24'h000000}, {10{24'h0}}};
					10'd25 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h545308}, {24'hfffd02}, {24'hfefd8f}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb1}, {24'hfffd52}, {24'hfffd00}, {24'he2ef5f}, {24'hc6e0dd}, {24'hf9fbb1}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'h82825c}, {24'h000000}, {10{24'h0}}};
					10'd26 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h848307}, {24'hfffd23}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfffd6f}, {24'hfffd06}, {24'hf6f91d}, {24'hc0dde4}, {24'hf9fab7}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfcfbb0}, {24'h424230}, {24'h000000}, {10{24'h0}}};
					10'd27 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'hadac0d}, {24'hfbfb84}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefd95}, {24'hfffd0b}, {24'hfefd03}, {24'hcde4a8}, {24'heaf3c6}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hafae7c}, {24'h060604}, {24'h000000}, {10{24'h0}}};
					10'd28 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h060602}, {24'hc7cd39}, {24'hd9ead4}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefda5}, {24'hfffd33}, {24'hfffd00}, {24'hfcfc23}, {24'he0eec5}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hd3d295}, {24'h1d1d15}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd29 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h242508}, {24'hc3d9a6}, {24'hcae2e7}, {24'hfefdb2}, {24'hfefdab}, {24'hfffd2f}, {24'hfffd00}, {24'hfffd29}, {24'hfefd9e}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hd0cf93}, {24'h12120d}, {24'h000000}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd30 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h858822}, {24'hbfdde2}, {24'hedf4c4}, {24'hfefdb1}, {24'hfefd62}, {24'hfffd03}, {24'hfffd10}, {24'hfefd95}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb1}, {24'hc5c48b}, {24'h222219}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					10'd31 : pattern <= {{24'h000000}, {24'h000000}, {24'h000000}, {24'h030404}, {24'hb0cbc2}, {24'hdaead6}, {24'hfefdb2}, {24'hfefd76}, {24'hfffd02}, {24'hfffd17}, {24'hfefd8b}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hfefdb2}, {24'hc0bf86}, {24'h161610}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {24'h000000}, {10{24'h0}}};
					default : pattern <= {32{24'h0}};
				endcase
			end
			default : begin
				pattern <= {32{24'h0}};
			end
		endcase
	end
endmodule
