/*
 * Avalon memory-mapped peripheral that generates VGA
 *
 * Stephen A. Edwards
 * Columbia University
 */

module vga_ball(input logic        	clk,
				input logic 	   	reset,
				input logic [31:0]  writedata,
				input logic 	   	write,
				input logic			chipselect,
				input logic [15:0]  address,

				output logic [7:0] 	VGA_R, VGA_G, VGA_B,
				output logic 	   	VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n,
				output logic 	   	VGA_SYNC_n);

	logic [10:0]	hcount;
	logic [9:0]     vcount;

	logic [7:0] 	color_r, color_g, color_b;
	logic [10:0]	x_cord;
	logic [9:0] 	y_cord;

	vga_counters counters(.clk50(clk), .*);

	always_ff @(posedge clk)
		if (reset) begin
			color_r <= 8'h80;
			color_g <= 8'h0;
			color_b <= 8'h80;
			x_cord <= 11'd1000;
			y_cord <= 10'd200;
			
		end else if (chipselect && write) begin
			case (address)
				// 3'h0 : x_cord <= writedata<<4;
				// 3'h1 : y_cord <= writedata<<3;
				3'h0 : color_r <= writedata[7:0];
				3'h1 : color_g <= writedata[7:0];
				3'h2 : color_b <= writedata[7:0];
				// x (0 - 639) or y (0 - 479) coords one at a time
				3'h3 : x_cord <= (writedata[10:0]<<1);
				3'h4 : y_cord <= (writedata[9:0]);
			endcase
		end
	always_comb begin
		{VGA_R, VGA_G, VGA_B} = {8'h10, 8'h20, 8'h30};
		// {x_cord, y_cord} = {11'd1000, 10'd231};
		if (VGA_BLANK_n)
			// if (((((hcount-x_cord)>>1)**2) + ((vcount-y_cord)**2)) <= 64)
			if (hcount > (x_cord-8) && hcount < (x_cord+8)) begin
				if ((vcount > (239) && vcount < (y_cord)))
					{VGA_R, VGA_G, VGA_B} = {8'hff, 8'hff, 8'hff};
				else if ((vcount < (239) && vcount > (y_cord)))
					{VGA_R, VGA_G, VGA_B} = {8'hff, 8'hff, 8'hff};
				else
					{VGA_R, VGA_G, VGA_B} = {color_r, color_g, color_b};
			end
			else
				{VGA_R, VGA_G, VGA_B} =
					{color_r, color_g, color_b};
	end

endmodule

module vga_counters(input logic 	     clk50, reset,
					output logic [10:0] hcount,  // hcount[10:1] is pixel column
					output logic [9:0]  vcount,  // vcount[9:0] is pixel row
					output logic 	     VGA_CLK, VGA_HS, VGA_VS, VGA_BLANK_n, VGA_SYNC_n);

/*
 * 640 X 480 VGA timing for a 50 MHz clock: one pixel every other cycle
 * 
 * HCOUNT 1599 0             1279       1599 0
 *             _______________              ________
 * ___________|    Video      |____________|  Video
 * 
 * 
 * |SYNC| BP |<-- HACTIVE -->|FP|SYNC| BP |<-- HACTIVE
 *       _______________________      _____________
 * |____|       VGA_HS          |____|
 */
// Parameters for hcount
	parameter 
		  HACTIVE      = 11'd 1280,
		  HFRONT_PORCH = 11'd 32,
		  HSYNC        = 11'd 192,
		  HBACK_PORCH  = 11'd 96,   
		  HTOTAL       = HACTIVE + HFRONT_PORCH + HSYNC +
		  HBACK_PORCH; // 1600

		  // Parameters for vcount
		  parameter 
		  VACTIVE      = 10'd 480,
		  VFRONT_PORCH = 10'd 10,
		  VSYNC        = 10'd 2,
		  VBACK_PORCH  = 10'd 33,
		  VTOTAL       = VACTIVE + VFRONT_PORCH + VSYNC +
		  VBACK_PORCH; // 525

		  logic endOfLine;

	always_ff @(posedge clk50 or posedge reset)
		if (reset)          hcount <= 0;
		else if (endOfLine) hcount <= 0;
		else  	         hcount <= hcount + 11'd 1;

	assign endOfLine = hcount == HTOTAL - 1;

	logic endOfField;

	always_ff @(posedge clk50 or posedge reset)
		if (reset)          vcount <= 0;
		else if (endOfLine)
			if (endOfField)   vcount <= 0;
			else              vcount <= vcount + 10'd 1;

	assign endOfField = vcount == VTOTAL - 1;

	// Horizontal sync: from 0x520 to 0x5DF (0x57F)
	// 101 0010 0000 to 101 1101 1111
	assign VGA_HS = !( (hcount[10:8] == 3'b101) &
					!(hcount[7:5] == 3'b111));
	assign VGA_VS = !( vcount[9:1] == (VACTIVE + VFRONT_PORCH) / 2);

	assign VGA_SYNC_n = 1'b0; // For putting sync on the green signal; unused

	// Horizontal active: 0 to 1279     Vertical active: 0 to 479
	// 101 0000 0000  1280	       01 1110 0000  480
	// 110 0011 1111  1599	       10 0000 1100  524
	assign VGA_BLANK_n = 	!( hcount[10] & (hcount[9] | hcount[8]) ) &
							!( vcount[9] | (vcount[8:5] == 4'b1111) );

		/* VGA_CLK is 25 MHz
		 *             __    __    __
		 * clk50    __|  |__|  |__|
		 *        
		 *             _____       __
		 * hcount[0]__|     |_____|
		 */
	assign VGA_CLK = hcount[0]; // 25 MHz clock: rising edge sensitive

endmodule
